module and_module(input wire a,b, output wire f);
    and(f,a,b);
endmodule
